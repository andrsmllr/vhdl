--============================================================================
--!
--! \file      <FILE_NAME>
--!
--! \project   <PROJECT_NAME>
--!
--! \langv     VHDL-2008
--!
--! \brief     <BRIEF_DESCRIPTION>.
--!
--! \details   <DETAILED_DESCRIPTION>.
--!
--! \bug       <BUGS_OR_KNOWN_ISSUES>.
--!
--! \see       <REFERENCES>
--!
--! \copyright <COPYRIGHT_OR_LICENSE>
--!
--! Revision history:
--!
--! \version   <VERSION>
--! \date      <YYYY-MM-DD>
--! \author    <AUTHOR_NAME>
--!
--============================================================================


library ieee;
    use ieee.numeric_std.all;
    use ieee.std_logic_1164.all;

package template_package is
end package template_package;

package body template_package is
end package body template_package;
