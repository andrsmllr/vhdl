--============================================================================
--!
--! \file      architecture_declaration.vhdl-2002.vhdl
--!
--! \project   vhdl_tutorial
--!
--! \langv     VHDL-2002
--!
--! \brief     Architecture declaration.
--!
--! \details   -
--!
--! \bug       -
--!
--! \see       "THE DESIGNER'S GUIDE TO VHDL THIRD EDITION", Peter J. Ashenden
--!
--! \copyright GPLv2
--!
--! Revision history:
--!
--! \version   1.0
--! \date      2015-12-29
--! \author    Andreas Muller
--!
--============================================================================

architecture architecture_vhdl_2002 of entity_vhdl_2002 is
begin
end architecture architecture_vhdl_2002;

