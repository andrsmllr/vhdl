--============================================================================
--!
--! \file      architecture_declaration.vhdl-1993.vhdl
--!
--! \project   vhdl_tutorial
--!
--! \langv     VHDL-1993
--!
--! \brief     Architecture declaration.
--!
--! \details   -
--!
--! \bug       -
--!
--! \see       "THE DESIGNER'S GUIDE TO VHDL THIRD EDITION", Peter J. Ashenden
--!
--! \copyright GPLv2
--!
--! Revision history:
--!
--! \version   1.0
--! \date      2015-12-29
--! \author    Andreas Muller
--!
--============================================================================

architecture architecture_vhdl_1993 of entity_vhdl_1993 is
begin
end architecture architecture_vhdl_1993;

