--============================================================================
--!
--! \file      mpeg2ts_pkg
--!
--! \project   mpeg2_lib
--!
--! \langv     VHDL-2002
--!
--! \brief     -
--!
--! \details   -
--!
--! \bug       -
--!
--! \see       -
--!
--! \copyright GPLv2
--!
--! Revision history:
--!
--! \version   0.1
--! \date      2015-06-06
--! \author    Andreas Mueller
--!
--============================================================================


library ieee;
    use ieee.numeric_std.all;
    use ieee.std_logic_1164.all;

package mpeg2ts_pkg is
end package mpeg2ts_pkg;

package body mpeg2ts_pkg is
end package body mpeg2ts_pkg;
