--============================================================================
--!
--! \file      component_declaration.vhdl-1987.vhdl
--!
--! \project   vhdl_tutorial
--!
--! \langv     VHDL-1987
--!
--! \brief     Component declaration.
--!
--! \details   -
--!
--! \bug       -
--!
--! \see       "THE DESIGNER'S GUIDE TO VHDL THIRD EDITION", Peter J. Ashenden
--!
--! \copyright GPLv2
--!
--! Revision history:
--!
--! \version   1.0
--! \date      2015-12-29
--! \author    Andreas Muller
--!
--============================================================================

component component_vhdl_1987
end component;

