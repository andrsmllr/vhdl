--============================================================================
--!
--! \file      architecture_declaration.vhdl-1987.vhdl
--!
--! \project   vhdl_tutorial
--!
--! \langv     VHDL-1987
--!
--! \brief     Architecture declaration.
--!
--! \details   -
--!
--! \bug       -
--!
--! \see       "THE DESIGNER'S GUIDE TO VHDL THIRD EDITION", Peter J. Ashenden
--!
--! \copyright GPLv2
--!
--! Revision history:
--!
--! \version   1.0
--! \date      2015-12-29
--! \author    Andreas Muller
--!
--============================================================================

architecture architecture_vhdl_1987 of entity_vhdl_1987 is
begin
end architecture_vhdl_1987;

