--============================================================================
--!
--! \file      entity_declaration.vhdl-1987.vhdl
--!
--! \project   vhdl_tutorial
--!
--! \langv     VHDL-1987
--!
--! \brief     Entity declaration.
--!
--! \details   -
--!
--! \bug       -
--!
--! \see       "THE DESIGNER'S GUIDE TO VHDL THIRD EDITION", Peter J. Ashenden
--!
--! \copyright GPLv2
--!
--! Revision history:
--!
--! \version   1.0
--! \date      2015-12-29
--! \author    Andreas Muller
--!
--============================================================================

entity entity_vhdl_1987 is
end entity_vhdl_1987;

